// --------------------------------------------------------------------
// >>>>>>>>>>>>>>>>>>>>>>>>> COPYRIGHT NOTICE <<<<<<<<<<<<<<<<<<<<<<<<<
// --------------------------------------------------------------------
// Module: LCD_RAM
// 
// Author: Step
// 
// Description: LCD_RAM
// 
// Web: www.stepfpga.com
//
// --------------------------------------------------------------------
// Code Revision History :
// --------------------------------------------------------------------
// Version: |Mod. Date:   |Changes Made:
// V1.1     |2016/10/30   |Initial ver
// --------------------------------------------------------------------
`timescale 1 ns / 100 ps
module LCD_RAM (Address, Q);

    input wire [7:0] Address;
    output reg [131:0] Q;
	 
	always @ (*)
		case(Address)
			8'd0  : Q = 132'h00000000000000000000000000000000;
			8'd1  : Q = 132'h00000000000000000000000000000000;
			8'd2  : Q = 132'h00000000000000000000000000000000;
			8'd3  : Q = 132'h00000000000000000000000000000000;
			8'd4  : Q = 132'h00000000000000000000000000000000;
			8'd5  : Q = 132'h00000000000000000000000000000000;
			8'd6  : Q = 132'h00000000000000000000000000000000;
			8'd7  : Q = 132'h00000000000000000000000000000000;
			8'd8  : Q = 132'h00000000000000000000000000000000;
			8'd9  : Q = 132'h00000000000000000000000000000000;
			8'd10 : Q = 132'h00000000000000000000000000000000;
			8'd11 : Q = 132'h00000000000000000000000000000000;
			8'd12 : Q = 132'h00000000000000000000000000000000;
			8'd13 : Q = 132'h00000000000000000000000000000000;
			8'd14 : Q = 132'h00000000000000000000000000000000;
			8'd15 : Q = 132'h00000000000000000000000000000000;
			8'd16 : Q = 132'h00000000000000000000000000000000;
			8'd17 : Q = 132'h00000000000000000000000000000000;
			8'd18 : Q = 132'h00000000000000000000000000000000;
			8'd19 : Q = 132'h00000000000000000000000000000000;
			8'd20 : Q = 132'h00000000000000000000000000000000;
			8'd21 : Q = 132'h00000000000000000000000000000000;
			8'd22 : Q = 132'h00000000000000000000000000000000;
			8'd23 : Q = 132'h00000000000000000000000000000000;
			8'd24 : Q = 132'h00000000000000000000000000000000;
			8'd25 : Q = 132'h00000000000000000000000000000000;
			8'd26 : Q = 132'h00000000000000000000000000000000;
			8'd27 : Q = 132'h00000000000000000000000000000000;
			8'd28 : Q = 132'h00000000000000000000000000000000;
			8'd29 : Q = 132'h00000000000000000000000000000000;
			8'd30 : Q = 132'h00000000000000000000000000000000;
			8'd31 : Q = 132'h00000000000000000000000000000000;
			8'd32 : Q = 132'h00000000000000FF8000000000000000;
			8'd33 : Q = 132'h00000000000003FFE000000000000000;
			8'd34 : Q = 132'h0000000000000FFFF800000000000000;
			8'd35 : Q = 132'h0000000000001FFFFC00000000000000;
			8'd36 : Q = 132'h0000000000003FFFFE00000000000000;
			8'd37 : Q = 132'h0000000000007FFFFF00000000000000;
			8'd38 : Q = 132'h000000000000FFFFFF80000000000000;
			8'd39 : Q = 132'h000000000000FFFFFF80000000000000;
			8'd40 : Q = 132'h000000000001FFFFFFC0000000000000;
			8'd41 : Q = 132'h000000000001FFFFFFC0000000000000;
			8'd42 : Q = 132'h000000000001FFC1FFC0000000000000;
			8'd43 : Q = 132'h000000000001FF80FFC0000000000000;
			8'd44 : Q = 132'h000000000001FF00FFC0000000000000;
			8'd45 : Q = 132'h000000000001FF007FC0000000000000;
			8'd46 : Q = 132'h000000000001FF00FFC0000000000000;
			8'd47 : Q = 132'h000000000001FF80FFC0000000000000;
			8'd48 : Q = 132'h000000000001FF81FFC0000000000000;
			8'd49 : Q = 132'h000000000001FFE3FFC0000000000000;
			8'd50 : Q = 132'h000000000001FFE7FFC0000000000000;
			8'd51 : Q = 132'h000000000000FFE7FF80000000000000;
			8'd52 : Q = 132'h000000000000FFE7FF80000007FC0000;
			8'd53 : Q = 132'h0000000000007FE7FF0000001FFF0000;
			8'd54 : Q = 132'h0000380000007FE7FE0000007FFF8000;
			8'd55 : Q = 132'h0001FF8000003FE7FC000000FFFFC000;
			8'd56 : Q = 132'h0007FFE000003FE7FC000001FFFFE000;
			8'd57 : Q = 132'h000FFFF000003FE7F8000003FFFFF000;
			8'd58 : Q = 132'h001FFFF800001FC7F8000003FFFFF000;
			8'd59 : Q = 132'h003FFFFC00001FC7F0000007FFFFF800;
			8'd60 : Q = 132'h003FFFFC00000FC7F0000007FFBFF800;
			8'd61 : Q = 132'h007FFFFE00000FCFF0000007FE0FFC00;
			8'd62 : Q = 132'h007F83FE00000FCFE000000FFC07FC00;
			8'd63 : Q = 132'h00FF01FE000007CFE000000FFC03FC00;
			8'd64 : Q = 132'h00FF00FE000007CFE000000FFC03FC00;
			8'd65 : Q = 132'h00FF00FE000007CFC000000FFC03FC00;
			8'd66 : Q = 132'h00FF00FE000007CFC000000FFC07FC00;
			8'd67 : Q = 132'h00FF01FE000007CFC000000FFC0FFC00;
			8'd68 : Q = 132'h007F81FE000007CFC000001FF81FF800;
			8'd69 : Q = 132'h007FE1FE000007CF8000001FF8FFF800;
			8'd70 : Q = 132'h007FF1FE0000078F8000001FF1FFF000;
			8'd71 : Q = 132'h003FF8FE0000078F8000001FE3FFF000;
			8'd72 : Q = 132'h003FF8FE0000078F8000003FC7FFE000;
			8'd73 : Q = 132'h001FFCFE0000079F8000003FCFFFC000;
			8'd74 : Q = 132'h000FFC7E0000079F0000003F8FFF8000;
			8'd75 : Q = 132'h0007FE7F0000079F0000007F1FFF0000;
			8'd76 : Q = 132'h0001FE3F0000079F0000007E3FFE0000;
			8'd77 : Q = 132'h0000FF3F0000079F000000FC7FFC0000;
			8'd78 : Q = 132'h00003F1F0000071F000000FCFFF80000;
			8'd79 : Q = 132'h00001F9F0000071F000001F8FFE00000;
			8'd80 : Q = 132'h00000F8F0000071F000001F1FFC00000;
			8'd81 : Q = 132'h000007CF0000071F000003E3FF800000;
			8'd82 : Q = 132'h000003C780000F3F000003C7FE000000;
			8'd83 : Q = 132'h000001E780000F3F0000078FFC000000;
			8'd84 : Q = 132'h000001E380000F3F80000F8FF0000000;
			8'd85 : Q = 132'h000000F3C0000F3F80000F1FE0000000;
			8'd86 : Q = 132'h00000071C0001E3FC0001E3FC0000000;
			8'd87 : Q = 132'h00000079C0003E3FC0003C7F80000000;
			8'd88 : Q = 132'h00000038E0003E3FE00078FF00000000;
			8'd89 : Q = 132'h0000003CF0007E1FF001F0FC00000000;
			8'd90 : Q = 132'h0000001C7C00FE1FFC07F1F800000000;
			8'd91 : Q = 132'h0000001E3E03FC1FFFFFE3F000000000;
			8'd92 : Q = 132'h0000000F3FFFFC8FFFFFC7E000000000;
			8'd93 : Q = 132'h0000000F1FFFF8CFFFFF0FC000000000;
			8'd94 : Q = 132'h0000000F8FFFF1C7FFFE1FC000000000;
			8'd95 : Q = 132'h00000007C3FFE1E3FFFC3F8000000000;
			8'd96 : Q = 132'h00000007E1FF83F1FFF07F0000000000;
			8'd97 : Q = 132'h00000003F0000FF83FC0FE0000000000;
			8'd98 : Q = 132'h00000003FC003FFC0003FC0000000000;
			8'd99 : Q = 132'h00000001FF00FFFF000FFC0000000000;
			8'd100: Q = 132'h00000001FFFFFFFFE07FF80000000000;
			8'd101: Q = 132'h00000000FFFFFFFFFFFFF80000000000;
			8'd102: Q = 132'h00000000FFFFFFFFFFFFF00000000000;
			8'd103: Q = 132'h000000007FFFFFFFFFFFE00000000000;
			8'd104: Q = 132'h000000007FFFFFFFFFFFE00000000000;
			8'd105: Q = 132'h000000007FFFFFFFFFFFC00000000000;
			8'd106: Q = 132'h000000003FFFFFFFFFFFC00000000000;
			8'd107: Q = 132'h000000003FFFFFFFFFFFC00000000000;
			8'd108: Q = 132'h000000003FFFFFFFFFFF800000000000;
			8'd109: Q = 132'h000000001FFFFFFFFFFF800000000000;
			8'd110: Q = 132'h000000001FFFFFFFFFFF000000000000;
			8'd111: Q = 132'h000000000FFFFFFFFFFF000000000000;
			8'd112: Q = 132'h000000000FFFFFFFFFFF000000000000;
			8'd113: Q = 132'h000000000FFFFFFFFFFE000000000000;
			8'd114: Q = 132'h0000000007FFFFFFFFFE000000000000;
			8'd115: Q = 132'h0000000007FFFFFFFFFC000000000000;
			8'd116: Q = 132'h0000000007FFFFFFFFFC000000000000;
			8'd117: Q = 132'h0000000003FFFFFFFFFC000000000000;
			8'd118: Q = 132'h0000000003FFFFFFFFF8000000000000;
			8'd119: Q = 132'h0000000003FFFFFFFFF8000000000000;
			8'd120: Q = 132'h0000000001FFFFFFFFF8000000000000;
			8'd121: Q = 132'h0000000001FFFFFFFFF0000000000000;
			8'd122: Q = 132'h0000000001FFFFFFFFF0000000000000;
			8'd123: Q = 132'h0000000000FFFFFFFFE0000000000000;
			8'd124: Q = 132'h0000000000FFFFFFFFE0000000000000;
			8'd125: Q = 132'h00000000007FFFFFFFC0000000000000;
			8'd126: Q = 132'h00000000003FFFFFFFC0000000000000;
			8'd127: Q = 132'h00000000003FFFFFFF80000000000000;
			8'd128: Q = 132'h00000000001FFFFFFF00000000000000;
			8'd129: Q = 132'h00000000000FFFFFFE00000000000000;
			8'd130: Q = 132'h000000000007FFFFFC00000000000000;
			8'd131: Q = 132'h000000000003FFFFF800000000000000;
			8'd132: Q = 132'h000000000000FFFFE000000000000000;
			8'd133: Q = 132'h0000000000001FFF8000000000000000;
			8'd134: Q = 132'h00000000000003F80000000000000000;
			8'd135: Q = 132'h00000000000000000000000000000000;
			8'd136: Q = 132'h00000000000000000000000000000000;
			8'd137: Q = 132'h00000000000000000000000000000000;
			8'd138: Q = 132'h00000000000000000000000000000000;
			8'd139: Q = 132'h00000000000000000000000000000000;
			8'd140: Q = 132'h00000000000000000000000000000000;
			8'd141: Q = 132'h00000000000000000000000000000000;
			8'd142: Q = 132'h00000000000000000000000000000000;
			8'd143: Q = 132'h00000000000000000000000000000000;
			8'd144: Q = 132'h00000000000000000000000000000000;
			8'd145: Q = 132'h00000000000000000000000000000000;
			8'd146: Q = 132'h00000000000000000000000000000000;
			8'd147: Q = 132'h00000000000000000000000000000000;
			8'd148: Q = 132'h00000000000000000000000000000000;
			8'd149: Q = 132'h00000000000000000000000000000000;
			8'd150: Q = 132'h00000000000000000000000000000000;
			8'd151: Q = 132'h00000000000000000000000000000000;
			8'd152: Q = 132'h00000000000000000000000000000000;
			8'd153: Q = 132'h00000000000000000000000000000000;
			8'd154: Q = 132'h00000000000000000000000000000000;
			8'd155: Q = 132'h00000000000000000000000000000000;
			8'd156: Q = 132'h00000000000000000000000000000000;
			8'd157: Q = 132'h00000000000000000000000000000000;
			8'd158: Q = 132'h00000000000000000000000000000000;
			8'd159: Q = 132'h00000000000000000000000000000000;
			default:Q = 132'h00000000000000000000000000000000;
		endcase
		
endmodule
