// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.9.0.99.2
// Netlist written on Thu Jan 24 14:52:31 2019
//
// Verilog Description of module Type_system
//

module Type_system (clk, rst_n, col, row, seg_1, seg_2) /* synthesis syn_module_defined=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(18[8:19])
    input clk;   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(20[11:14])
    input rst_n;   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(21[11:16])
    input [3:0]col;   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(22[15:18])
    output [3:0]row;   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(23[16:19])
    output [8:0]seg_1;   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(24[16:21])
    output [8:0]seg_2;   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(25[16:21])
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(20[11:14])
    
    wire rst_n_c, col_c_3, col_c_2, col_c_1, col_c_0, row_c_3, row_c_2, 
        row_c_1, row_c_0, seg_1_c_5, seg_2_c_6, seg_2_c_5, seg_2_c_4, 
        seg_2_c_3, seg_2_c_2, seg_2_c_1, seg_2_c_0;
    wire [15:0]key_pulse;   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(29[15:24])
    wire [7:0]seg_data;   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(41[14:22])
    
    wire VCC_net;
    wire [15:0]key_out_adj_154;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(27[20:27])
    wire [15:0]cnt;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(44[15:18])
    wire [15:0]key_out_r;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(97[15:24])
    
    wire rst_n_N_6, GND_net, n1032, n5;
    
    VHI i5 (.Z(VCC_net));
    OB row_pad_3 (.I(row_c_3), .O(row[3]));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(23[16:19])
    VLO i1 (.Z(GND_net));
    TSALL TSALL_INST (.TSALL(GND_net));
    Decoder u2 (.\key_out_r[15] (key_out_r[15]), .\key_out[15] (key_out_adj_154[15]), 
            .key_pulse({key_pulse}), .\key_out_r[0] (key_out_r[0]), .\key_out[0] (key_out_adj_154[0]), 
            .\key_out_r[1] (key_out_r[1]), .\key_out[1] (key_out_adj_154[1]), 
            .\key_out_r[6] (key_out_r[6]), .\key_out[6] (key_out_adj_154[6]), 
            .\key_out_r[7] (key_out_r[7]), .\key_out[7] (key_out_adj_154[7]), 
            .\key_out_r[4] (key_out_r[4]), .\key_out[4] (key_out_adj_154[4]), 
            .\key_out_r[5] (key_out_r[5]), .\key_out[5] (key_out_adj_154[5]), 
            .rst_n_c(rst_n_c), .rst_n_N_6(rst_n_N_6), .\seg_data[4] (seg_data[4]), 
            .clk_c(clk_c), .\key_out_r[9] (key_out_r[9]), .\key_out[9] (key_out_adj_154[9]), 
            .\seg_data[3] (seg_data[3]), .\seg_data[2] (seg_data[2]), .\seg_data[1] (seg_data[1]), 
            .\key_out_r[13] (key_out_r[13]), .\key_out[13] (key_out_adj_154[13]), 
            .\seg_data[0] (seg_data[0]), .\key_out_r[11] (key_out_r[11]), 
            .\key_out[11] (key_out_adj_154[11])) /* synthesis syn_module_defined=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(43[9] 49[2])
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    IB col_pad_0 (.I(col[0]), .O(col_c_0));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(22[15:18])
    IB col_pad_1 (.I(col[1]), .O(col_c_1));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(22[15:18])
    IB col_pad_2 (.I(col[2]), .O(col_c_2));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(22[15:18])
    IB col_pad_3 (.I(col[3]), .O(col_c_3));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(22[15:18])
    IB rst_n_pad (.I(rst_n), .O(rst_n_c));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(21[11:16])
    IB clk_pad (.I(clk), .O(clk_c));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(20[11:14])
    OB seg_2_pad_0 (.I(seg_2_c_0), .O(seg_2[0]));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(25[16:21])
    OB seg_2_pad_1 (.I(seg_2_c_1), .O(seg_2[1]));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(25[16:21])
    OB seg_2_pad_2 (.I(seg_2_c_2), .O(seg_2[2]));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(25[16:21])
    OB seg_2_pad_3 (.I(seg_2_c_3), .O(seg_2[3]));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(25[16:21])
    OB seg_2_pad_4 (.I(seg_2_c_4), .O(seg_2[4]));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(25[16:21])
    OB seg_2_pad_5 (.I(seg_2_c_5), .O(seg_2[5]));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(25[16:21])
    OB seg_2_pad_6 (.I(seg_2_c_6), .O(seg_2[6]));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(25[16:21])
    OB seg_2_pad_7 (.I(GND_net), .O(seg_2[7]));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(25[16:21])
    OB seg_2_pad_8 (.I(GND_net), .O(seg_2[8]));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(25[16:21])
    OB seg_1_pad_0 (.I(seg_1_c_5), .O(seg_1[0]));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(24[16:21])
    OB seg_1_pad_1 (.I(VCC_net), .O(seg_1[1]));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(24[16:21])
    OB seg_1_pad_2 (.I(VCC_net), .O(seg_1[2]));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(24[16:21])
    OB seg_1_pad_3 (.I(seg_1_c_5), .O(seg_1[3]));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(24[16:21])
    OB seg_1_pad_4 (.I(seg_1_c_5), .O(seg_1[4]));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(24[16:21])
    OB seg_1_pad_5 (.I(seg_1_c_5), .O(seg_1[5]));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(24[16:21])
    OB seg_1_pad_6 (.I(GND_net), .O(seg_1[6]));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(24[16:21])
    OB seg_1_pad_7 (.I(GND_net), .O(seg_1[7]));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(24[16:21])
    OB seg_1_pad_8 (.I(GND_net), .O(seg_1[8]));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(24[16:21])
    OB row_pad_0 (.I(row_c_0), .O(row[0]));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(23[16:19])
    OB row_pad_1 (.I(row_c_1), .O(row[1]));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(23[16:19])
    OB row_pad_2 (.I(row_c_2), .O(row[2]));   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(23[16:19])
    LUT4 i682_2_lut_3_lut_4_lut (.A(cnt[0]), .B(n5), .C(cnt[13]), .D(cnt[12]), 
         .Z(n1032)) /* synthesis lut_function=(!((B (C (D)))+!A)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(55[12:22])
    defparam i682_2_lut_3_lut_4_lut.init = 16'h2aaa;
    GSR GSR_INST (.GSR(VCC_net));
    Segment_led u4 (.\seg_data[0] (seg_data[0]), .\seg_data[2] (seg_data[2]), 
            .\seg_data[3] (seg_data[3]), .\seg_data[1] (seg_data[1]), .seg_2_c_0(seg_2_c_0), 
            .seg_2_c_5(seg_2_c_5), .seg_2_c_6(seg_2_c_6), .seg_2_c_1(seg_2_c_1), 
            .seg_2_c_4(seg_2_c_4), .seg_2_c_2(seg_2_c_2), .seg_2_c_3(seg_2_c_3)) /* synthesis syn_module_defined=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(59[13] 63[2])
    Segment_led_U0 u3 (.\seg_data[4] (seg_data[4]), .seg_1_c_5(seg_1_c_5)) /* synthesis syn_module_defined=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(52[13] 56[2])
    Array_KeyBoard u1 (.clk_c(clk_c), .rst_n_N_6(rst_n_N_6), .key_pulse({key_pulse}), 
            .\key_out[9] (key_out_adj_154[9]), .\key_out_r[13] (key_out_r[13]), 
            .\key_out[13] (key_out_adj_154[13]), .col_c_1(col_c_1), .col_c_0(col_c_0), 
            .\key_out_r[0] (key_out_r[0]), .\key_out[0] (key_out_adj_154[0]), 
            .\cnt[0] (cnt[0]), .n5(n5), .\cnt[13] (cnt[13]), .\cnt[12] (cnt[12]), 
            .\key_out[7] (key_out_adj_154[7]), .\key_out_r[9] (key_out_r[9]), 
            .\key_out[6] (key_out_adj_154[6]), .\key_out_r[11] (key_out_r[11]), 
            .\key_out[11] (key_out_adj_154[11]), .\key_out[5] (key_out_adj_154[5]), 
            .\key_out[4] (key_out_adj_154[4]), .\key_out_r[1] (key_out_r[1]), 
            .\key_out[1] (key_out_adj_154[1]), .\key_out_r[4] (key_out_r[4]), 
            .\key_out_r[15] (key_out_r[15]), .\key_out[15] (key_out_adj_154[15]), 
            .\key_out_r[5] (key_out_r[5]), .GND_net(GND_net), .row_c_2(row_c_2), 
            .VCC_net(VCC_net), .row_c_1(row_c_1), .row_c_0(row_c_0), .n1032(n1032), 
            .\key_out_r[7] (key_out_r[7]), .\key_out_r[6] (key_out_r[6]), 
            .col_c_3(col_c_3), .col_c_2(col_c_2), .row_c_3(row_c_3)) /* synthesis syn_module_defined=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(31[16] 39[2])
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module Decoder
//

module Decoder (\key_out_r[15] , \key_out[15] , key_pulse, \key_out_r[0] , 
            \key_out[0] , \key_out_r[1] , \key_out[1] , \key_out_r[6] , 
            \key_out[6] , \key_out_r[7] , \key_out[7] , \key_out_r[4] , 
            \key_out[4] , \key_out_r[5] , \key_out[5] , rst_n_c, rst_n_N_6, 
            \seg_data[4] , clk_c, \key_out_r[9] , \key_out[9] , \seg_data[3] , 
            \seg_data[2] , \seg_data[1] , \key_out_r[13] , \key_out[13] , 
            \seg_data[0] , \key_out_r[11] , \key_out[11] ) /* synthesis syn_module_defined=1 */ ;
    input \key_out_r[15] ;
    input \key_out[15] ;
    input [15:0]key_pulse;
    input \key_out_r[0] ;
    input \key_out[0] ;
    input \key_out_r[1] ;
    input \key_out[1] ;
    input \key_out_r[6] ;
    input \key_out[6] ;
    input \key_out_r[7] ;
    input \key_out[7] ;
    input \key_out_r[4] ;
    input \key_out[4] ;
    input \key_out_r[5] ;
    input \key_out[5] ;
    input rst_n_c;
    output rst_n_N_6;
    output \seg_data[4] ;
    input clk_c;
    input \key_out_r[9] ;
    input \key_out[9] ;
    output \seg_data[3] ;
    output \seg_data[2] ;
    output \seg_data[1] ;
    input \key_out_r[13] ;
    input \key_out[13] ;
    output \seg_data[0] ;
    input \key_out_r[11] ;
    input \key_out[11] ;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(20[11:14])
    
    wire n709, n686, n812, n756, n1044, n707, n17, n687, n704, 
        n21, n20, n670, n702, n676, n1042, n6, n653, n705, 
        n770, n668, n681, n1167, n703, n1153, n706, n675, n662, 
        n748, n1045, n26, n19, n29, n4, n1179, clk_c_enable_5, 
        n1158, n684, n708, n663, n746, n698, n32;
    
    LUT4 i844_4_lut (.A(n709), .B(n686), .C(n812), .D(n756), .Z(n1044)) /* synthesis lut_function=(!(A (B (C (D))))) */ ;
    defparam i844_4_lut.init = 16'h7fff;
    LUT4 i2_3_lut_4_lut (.A(\key_out_r[15] ), .B(\key_out[15] ), .C(n707), 
         .D(key_pulse[14]), .Z(n709)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (C+!(D))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(46[4:12])
    defparam i2_3_lut_4_lut.init = 16'hf2ff;
    LUT4 key_pulse_15__I_0_40_i17_2_lut_4_lut (.A(\key_out_r[0] ), .B(\key_out[0] ), 
         .C(\key_out_r[1] ), .D(\key_out[1] ), .Z(n17)) /* synthesis lut_function=(!(A (B ((D)+!C))+!A ((D)+!C))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(46[4:12])
    defparam key_pulse_15__I_0_40_i17_2_lut_4_lut.init = 16'h22f2;
    LUT4 i1_2_lut_3_lut (.A(key_pulse[12]), .B(key_pulse[13]), .C(n687), 
         .Z(n707)) /* synthesis lut_function=(A+(B+(C))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(42[4:12])
    defparam i1_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_adj_3 (.A(key_pulse[14]), .B(key_pulse[15]), .C(n687), 
         .Z(n704)) /* synthesis lut_function=(A+(B+(C))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(45[4:12])
    defparam i1_2_lut_3_lut_adj_3.init = 16'hfefe;
    LUT4 key_pulse_15__I_0_40_i21_2_lut_4_lut (.A(\key_out_r[6] ), .B(\key_out[6] ), 
         .C(\key_out_r[7] ), .D(\key_out[7] ), .Z(n21)) /* synthesis lut_function=(!(A (B ((D)+!C))+!A ((D)+!C))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(46[4:12])
    defparam key_pulse_15__I_0_40_i21_2_lut_4_lut.init = 16'h22f2;
    LUT4 key_pulse_15__I_0_40_i20_2_lut_4_lut (.A(\key_out_r[4] ), .B(\key_out[4] ), 
         .C(\key_out_r[5] ), .D(\key_out[5] ), .Z(n20)) /* synthesis lut_function=(!(A (B ((D)+!C))+!A ((D)+!C))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(46[4:12])
    defparam key_pulse_15__I_0_40_i20_2_lut_4_lut.init = 16'h22f2;
    LUT4 i2_3_lut_4_lut_adj_4 (.A(n17), .B(n670), .C(key_pulse[2]), .D(key_pulse[3]), 
         .Z(n702)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(34[4:12])
    defparam i2_3_lut_4_lut_adj_4.init = 16'hffef;
    LUT4 i4_4_lut (.A(n676), .B(n686), .C(n1042), .D(n6), .Z(n653)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i4_4_lut.init = 16'hfff7;
    LUT4 i461_2_lut (.A(n705), .B(n770), .Z(n812)) /* synthesis lut_function=(A (B)) */ ;
    defparam i461_2_lut.init = 16'h8888;
    LUT4 i2_4_lut (.A(n668), .B(n681), .C(n1167), .D(n703), .Z(n1153)) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;
    defparam i2_4_lut.init = 16'hdfff;
    LUT4 i407_4_lut (.A(n706), .B(key_pulse[9]), .C(n675), .D(key_pulse[8]), 
         .Z(n756)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;
    defparam i407_4_lut.init = 16'haaa2;
    LUT4 i854_4_lut (.A(n662), .B(n702), .C(n812), .D(n748), .Z(n1045)) /* synthesis lut_function=(!(A (B (C (D))))) */ ;
    defparam i854_4_lut.init = 16'h7fff;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n20), .B(n21), .C(n26), .D(n19), .Z(n687)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(34[4:12])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_5 (.A(n20), .B(n21), .C(n29), .D(n26), 
         .Z(n670)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(34[4:12])
    defparam i1_2_lut_3_lut_4_lut_adj_5.init = 16'hfffe;
    LUT4 i2_3_lut_4_lut_adj_6 (.A(n17), .B(n670), .C(key_pulse[2]), .D(key_pulse[3]), 
         .Z(n703)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(34[4:12])
    defparam i2_3_lut_4_lut_adj_6.init = 16'hfeff;
    LUT4 i2_4_lut_adj_7 (.A(key_pulse[5]), .B(n21), .C(key_pulse[4]), 
         .D(n4), .Z(n668)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(37[4:12])
    defparam i2_4_lut_adj_7.init = 16'hfffd;
    LUT4 rst_n_I_0_1_lut (.A(rst_n_c), .Z(rst_n_N_6)) /* synthesis lut_function=(!(A)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(64[6:12])
    defparam rst_n_I_0_1_lut.init = 16'h5555;
    LUT4 i2_3_lut (.A(n1179), .B(n653), .C(n703), .Z(clk_c_enable_5)) /* synthesis lut_function=((B+!(C))+!A) */ ;
    defparam i2_3_lut.init = 16'hdfdf;
    LUT4 i1_2_lut_3_lut_adj_8 (.A(key_pulse[8]), .B(key_pulse[9]), .C(n1158), 
         .Z(n684)) /* synthesis lut_function=(A+(B+(C))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(46[4:12])
    defparam i1_2_lut_3_lut_adj_8.init = 16'hfefe;
    LUT4 i808_2_lut_4_lut (.A(key_pulse[13]), .B(n704), .C(key_pulse[12]), 
         .D(n708), .Z(n1167)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;
    defparam i808_2_lut_4_lut.init = 16'hfd00;
    FD1P3DX seg_data_i0_i4 (.D(n1044), .SP(clk_c_enable_5), .CK(clk_c), 
            .CD(rst_n_N_6), .Q(\seg_data[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=43, LSE_RLINE=49 */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(30[11] 50[5])
    defparam seg_data_i0_i4.GSR = "ENABLED";
    LUT4 i820_4_lut (.A(n756), .B(n770), .C(n663), .D(n748), .Z(n1179)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i820_4_lut.init = 16'h8000;
    LUT4 i841_2_lut_4_lut (.A(key_pulse[9]), .B(n675), .C(key_pulse[8]), 
         .D(n663), .Z(n746)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !(C+!(D))))) */ ;
    defparam i841_2_lut_4_lut.init = 16'h10ff;
    LUT4 i2_3_lut_4_lut_adj_9 (.A(\key_out_r[9] ), .B(\key_out[9] ), .C(n675), 
         .D(key_pulse[8]), .Z(n676)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (C+!(D))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(40[4:12])
    defparam i2_3_lut_4_lut_adj_9.init = 16'hf2ff;
    LUT4 i2_3_lut_4_lut_adj_10 (.A(n20), .B(n4), .C(key_pulse[6]), .D(key_pulse[7]), 
         .Z(n663)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(38[4:12])
    defparam i2_3_lut_4_lut_adj_10.init = 16'hfeff;
    LUT4 i2_3_lut_4_lut_adj_11 (.A(n20), .B(n4), .C(key_pulse[6]), .D(key_pulse[7]), 
         .Z(n662)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(38[4:12])
    defparam i2_3_lut_4_lut_adj_11.init = 16'hffef;
    LUT4 i1_2_lut_3_lut_adj_12 (.A(n26), .B(n29), .C(n19), .Z(n4)) /* synthesis lut_function=(A+(B+(C))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(32[4:12])
    defparam i1_2_lut_3_lut_adj_12.init = 16'hfefe;
    LUT4 i421_4_lut (.A(n708), .B(key_pulse[11]), .C(n684), .D(key_pulse[10]), 
         .Z(n770)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;
    defparam i421_4_lut.init = 16'haaa2;
    FD1P3DX seg_data_i0_i3 (.D(n746), .SP(clk_c_enable_5), .CK(clk_c), 
            .CD(rst_n_N_6), .Q(\seg_data[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=43, LSE_RLINE=49 */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(30[11] 50[5])
    defparam seg_data_i0_i3.GSR = "ENABLED";
    FD1P3DX seg_data_i0_i2 (.D(n1153), .SP(clk_c_enable_5), .CK(clk_c), 
            .CD(rst_n_N_6), .Q(\seg_data[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=43, LSE_RLINE=49 */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(30[11] 50[5])
    defparam seg_data_i0_i2.GSR = "ENABLED";
    FD1P3DX seg_data_i0_i1 (.D(n1045), .SP(clk_c_enable_5), .CK(clk_c), 
            .CD(rst_n_N_6), .Q(\seg_data[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=43, LSE_RLINE=49 */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(30[11] 50[5])
    defparam seg_data_i0_i1.GSR = "ENABLED";
    LUT4 i1_3_lut (.A(n681), .B(n702), .C(n705), .Z(n6)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i1_3_lut.init = 16'hbfbf;
    LUT4 i2_3_lut_4_lut_adj_13 (.A(\key_out_r[1] ), .B(\key_out[1] ), .C(n698), 
         .D(key_pulse[0]), .Z(n1042)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;
    defparam i2_3_lut_4_lut_adj_13.init = 16'h0d00;
    LUT4 i1_4_lut (.A(n709), .B(n32), .C(n4), .D(key_pulse[5]), .Z(n681)) /* synthesis lut_function=(!(A ((C+(D))+!B))) */ ;
    defparam i1_4_lut.init = 16'h555d;
    LUT4 i1_2_lut_3_lut_adj_14 (.A(key_pulse[10]), .B(key_pulse[11]), .C(n1158), 
         .Z(n675)) /* synthesis lut_function=(A+(B+(C))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(46[4:12])
    defparam i1_2_lut_3_lut_adj_14.init = 16'hfefe;
    LUT4 i1_4_lut_adj_15 (.A(\key_out_r[7] ), .B(key_pulse[6]), .C(\key_out[7] ), 
         .D(key_pulse[4]), .Z(n32)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C (D)))+!A (B (D)+!B !(D)))) */ ;
    defparam i1_4_lut_adj_15.init = 16'h31c4;
    LUT4 key_pulse_15__I_0_28_i26_2_lut_3_lut_4_lut (.A(key_pulse[10]), .B(key_pulse[11]), 
         .C(key_pulse[9]), .D(key_pulse[8]), .Z(n26)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(46[4:12])
    defparam key_pulse_15__I_0_28_i26_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 key_pulse_15__I_0_30_i19_2_lut_3_lut (.A(key_pulse[2]), .B(key_pulse[3]), 
         .C(n17), .Z(n19)) /* synthesis lut_function=(A+(B+(C))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(46[4:12])
    defparam key_pulse_15__I_0_30_i19_2_lut_3_lut.init = 16'hfefe;
    LUT4 i2_3_lut_4_lut_adj_16 (.A(\key_out_r[15] ), .B(\key_out[15] ), 
         .C(n707), .D(key_pulse[14]), .Z(n708)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(47[4:12])
    defparam i2_3_lut_4_lut_adj_16.init = 16'hfffd;
    LUT4 i1_2_lut_3_lut_adj_17 (.A(key_pulse[2]), .B(key_pulse[3]), .C(n670), 
         .Z(n698)) /* synthesis lut_function=(A+(B+(C))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(46[4:12])
    defparam i1_2_lut_3_lut_adj_17.init = 16'hfefe;
    LUT4 i2_3_lut_4_lut_adj_18 (.A(\key_out_r[13] ), .B(\key_out[13] ), 
         .C(n704), .D(key_pulse[12]), .Z(n705)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (C+!(D))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(44[4:12])
    defparam i2_3_lut_4_lut_adj_18.init = 16'hf2ff;
    LUT4 i1_2_lut_3_lut_4_lut_adj_19 (.A(n20), .B(n21), .C(n29), .D(n19), 
         .Z(n1158)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(34[4:12])
    defparam i1_2_lut_3_lut_4_lut_adj_19.init = 16'hfffe;
    LUT4 key_pulse_15__I_0_26_i29_2_lut_3_lut_4_lut (.A(key_pulse[12]), .B(key_pulse[13]), 
         .C(key_pulse[15]), .D(key_pulse[14]), .Z(n29)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(42[4:12])
    defparam key_pulse_15__I_0_26_i29_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_4_lut_adj_20 (.A(\key_out_r[13] ), .B(\key_out[13] ), 
         .C(n704), .D(key_pulse[12]), .Z(n706)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(45[4:12])
    defparam i2_3_lut_4_lut_adj_20.init = 16'hfffd;
    FD1P3DX seg_data_i0_i0 (.D(n653), .SP(clk_c_enable_5), .CK(clk_c), 
            .CD(rst_n_N_6), .Q(\seg_data[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=43, LSE_RLINE=49 */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(30[11] 50[5])
    defparam seg_data_i0_i0.GSR = "ENABLED";
    LUT4 i2_3_lut_4_lut_adj_21 (.A(\key_out_r[11] ), .B(\key_out[11] ), 
         .C(n684), .D(key_pulse[10]), .Z(n686)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (C+!(D))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/decoder.v(42[4:12])
    defparam i2_3_lut_4_lut_adj_21.init = 16'hf2ff;
    LUT4 i399_4_lut (.A(n668), .B(key_pulse[1]), .C(n698), .D(key_pulse[0]), 
         .Z(n748)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;
    defparam i399_4_lut.init = 16'haaa2;
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module Segment_led
//

module Segment_led (\seg_data[0] , \seg_data[2] , \seg_data[3] , \seg_data[1] , 
            seg_2_c_0, seg_2_c_5, seg_2_c_6, seg_2_c_1, seg_2_c_4, 
            seg_2_c_2, seg_2_c_3) /* synthesis syn_module_defined=1 */ ;
    input \seg_data[0] ;
    input \seg_data[2] ;
    input \seg_data[3] ;
    input \seg_data[1] ;
    output seg_2_c_0;
    output seg_2_c_5;
    output seg_2_c_6;
    output seg_2_c_1;
    output seg_2_c_4;
    output seg_2_c_2;
    output seg_2_c_3;
    
    
    LUT4 seg_data_3__I_0_Mux_0_i15_4_lut (.A(\seg_data[0] ), .B(\seg_data[2] ), 
         .C(\seg_data[3] ), .D(\seg_data[1] ), .Z(seg_2_c_0)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B (C (D))))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/segment_led.v(25[2] 37[9])
    defparam seg_data_3__I_0_Mux_0_i15_4_lut.init = 16'h0f39;
    LUT4 seg_data_0__bdd_4_lut_861 (.A(\seg_data[0] ), .B(\seg_data[3] ), 
         .C(\seg_data[2] ), .D(\seg_data[1] ), .Z(seg_2_c_5)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A (B (C+(D))+!B !(C+!(D))))) */ ;
    defparam seg_data_0__bdd_4_lut_861.init = 16'h103d;
    LUT4 seg_data_1__bdd_4_lut (.A(\seg_data[1] ), .B(\seg_data[0] ), .C(\seg_data[3] ), 
         .D(\seg_data[2] ), .Z(seg_2_c_6)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C))+!A (C (D)+!C !(D)))) */ ;
    defparam seg_data_1__bdd_4_lut.init = 16'h075a;
    LUT4 seg_data_0__bdd_4_lut_860 (.A(\seg_data[0] ), .B(\seg_data[3] ), 
         .C(\seg_data[2] ), .D(\seg_data[1] ), .Z(seg_2_c_1)) /* synthesis lut_function=(!(A (B (C+(D))+!B !((D)+!C))+!A (B (C+(D))+!B (C (D))))) */ ;
    defparam seg_data_0__bdd_4_lut_860.init = 16'h231f;
    LUT4 i847_4_lut (.A(\seg_data[0] ), .B(\seg_data[2] ), .C(\seg_data[3] ), 
         .D(\seg_data[1] ), .Z(seg_2_c_4)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B (C (D))))) */ ;
    defparam i847_4_lut.init = 16'h0511;
    LUT4 seg_data_1__bdd_4_lut_859 (.A(\seg_data[1] ), .B(\seg_data[0] ), 
         .C(\seg_data[3] ), .D(\seg_data[2] ), .Z(seg_2_c_2)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (C (D)))) */ ;
    defparam seg_data_1__bdd_4_lut_859.init = 16'h0f5d;
    LUT4 seg_data_0__bdd_4_lut (.A(\seg_data[0] ), .B(\seg_data[3] ), .C(\seg_data[1] ), 
         .D(\seg_data[2] ), .Z(seg_2_c_3)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C (D)+!C !(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;
    defparam seg_data_0__bdd_4_lut.init = 16'h123d;
    
endmodule
//
// Verilog Description of module Segment_led_U0
//

module Segment_led_U0 (\seg_data[4] , seg_1_c_5) /* synthesis syn_module_defined=1 */ ;
    input \seg_data[4] ;
    output seg_1_c_5;
    
    
    LUT4 i93_1_lut (.A(\seg_data[4] ), .Z(seg_1_c_5)) /* synthesis lut_function=(!(A)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/segment_led.v(25[2] 37[9])
    defparam i93_1_lut.init = 16'h5555;
    
endmodule
//
// Verilog Description of module Array_KeyBoard
//

module Array_KeyBoard (clk_c, rst_n_N_6, key_pulse, \key_out[9] , \key_out_r[13] , 
            \key_out[13] , col_c_1, col_c_0, \key_out_r[0] , \key_out[0] , 
            \cnt[0] , n5, \cnt[13] , \cnt[12] , \key_out[7] , \key_out_r[9] , 
            \key_out[6] , \key_out_r[11] , \key_out[11] , \key_out[5] , 
            \key_out[4] , \key_out_r[1] , \key_out[1] , \key_out_r[4] , 
            \key_out_r[15] , \key_out[15] , \key_out_r[5] , GND_net, 
            row_c_2, VCC_net, row_c_1, row_c_0, n1032, \key_out_r[7] , 
            \key_out_r[6] , col_c_3, col_c_2, row_c_3) /* synthesis syn_module_defined=1 */ ;
    input clk_c;
    input rst_n_N_6;
    output [15:0]key_pulse;
    output \key_out[9] ;
    output \key_out_r[13] ;
    output \key_out[13] ;
    input col_c_1;
    input col_c_0;
    output \key_out_r[0] ;
    output \key_out[0] ;
    output \cnt[0] ;
    output n5;
    output \cnt[13] ;
    output \cnt[12] ;
    output \key_out[7] ;
    output \key_out_r[9] ;
    output \key_out[6] ;
    output \key_out_r[11] ;
    output \key_out[11] ;
    output \key_out[5] ;
    output \key_out[4] ;
    output \key_out_r[1] ;
    output \key_out[1] ;
    output \key_out_r[4] ;
    output \key_out_r[15] ;
    output \key_out[15] ;
    output \key_out_r[5] ;
    input GND_net;
    output row_c_2;
    input VCC_net;
    output row_c_1;
    output row_c_0;
    input n1032;
    output \key_out_r[7] ;
    output \key_out_r[6] ;
    input col_c_3;
    input col_c_2;
    output row_c_3;
    
    wire clk_200hz_N_24 /* synthesis is_inv_clock=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(27[20:27])
    wire clk_200hz /* synthesis is_clock=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(45[10:19])
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/type_system.v(20[11:14])
    
    wire clk_200hz_N_25;
    wire [15:0]key_out_r;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(97[15:24])
    wire [15:0]key_out;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(27[20:27])
    
    wire clk_200hz_N_24_enable_45;
    wire [3:0]key_out_15__N_113;
    wire [15:0]key_r;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(79[17:22])
    
    wire clk_200hz_N_24_enable_48;
    wire [15:0]key;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(79[13:16])
    wire [3:0]key_out_15__N_117;
    wire [3:0]n68;
    wire [3:0]key_out_15__N_121;
    wire [14:0]n82;
    
    wire clk_200hz_N_24_enable_46, clk_200hz_N_26;
    wire [3:0]row_3__N_1;
    
    wire n20;
    wire [15:0]cnt;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(44[15:18])
    
    wire n4, n1047, n6, n1040, n1039, n1038, n1037, n1036, n1035, 
        n1034;
    wire [3:0]key_out_15__N_109;
    
    INV i900 (.A(clk_200hz), .Z(clk_200hz_N_24));
    FD1S3DX clk_200hz_38 (.D(clk_200hz_N_25), .CK(clk_c), .CD(rst_n_N_6), 
            .Q(clk_200hz)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(50[12] 58[6])
    defparam clk_200hz_38.GSR = "ENABLED";
    LUT4 key_out_r_15__I_0_i13_2_lut (.A(key_out_r[12]), .B(key_out[12]), 
         .Z(key_pulse[12])) /* synthesis lut_function=(!((B)+!A)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(105[20:43])
    defparam key_out_r_15__I_0_i13_2_lut.init = 16'h2222;
    FD1P3BX key_out_i9 (.D(key_out_15__N_113[1]), .SP(clk_200hz_N_24_enable_45), 
            .CK(clk_200hz_N_24), .PD(rst_n_N_6), .Q(\key_out[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_out_i9.GSR = "ENABLED";
    LUT4 key_out_r_15__I_0_i14_2_lut (.A(\key_out_r[13] ), .B(\key_out[13] ), 
         .Z(key_pulse[13])) /* synthesis lut_function=(!((B)+!A)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(105[20:43])
    defparam key_out_r_15__I_0_i14_2_lut.init = 16'h2222;
    FD1P3BX key_out_i8 (.D(key_out_15__N_113[0]), .SP(clk_200hz_N_24_enable_45), 
            .CK(clk_200hz_N_24), .PD(rst_n_N_6), .Q(key_out[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_out_i8.GSR = "ENABLED";
    FD1P3BX key_r_i0 (.D(key[0]), .SP(clk_200hz_N_24_enable_48), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key_r[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_r_i0.GSR = "ENABLED";
    FD1P3BX key_i1 (.D(col_c_1), .SP(clk_200hz_N_24_enable_48), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_i1.GSR = "ENABLED";
    FD1P3BX key_i0 (.D(col_c_0), .SP(clk_200hz_N_24_enable_48), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_i0.GSR = "ENABLED";
    LUT4 or_22_i4_2_lut (.A(key_r[7]), .B(key[7]), .Z(key_out_15__N_117[3])) /* synthesis lut_function=(A+(B)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(89[37:60])
    defparam or_22_i4_2_lut.init = 16'heeee;
    FD1S3BX key_out_r_i0 (.D(\key_out[0] ), .CK(clk_c), .PD(rst_n_N_6), 
            .Q(\key_out_r[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(101[9:30])
    defparam key_out_r_i0.GSR = "ENABLED";
    FD1P3BX key_r_i15 (.D(key[15]), .SP(n68[3]), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key_r[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_r_i15.GSR = "ENABLED";
    FD1P3BX key_out_i0 (.D(key_out_15__N_121[0]), .SP(clk_200hz_N_24_enable_48), 
            .CK(clk_200hz_N_24), .PD(rst_n_N_6), .Q(\key_out[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_out_i0.GSR = "ENABLED";
    FD1P3BX key_r_i14 (.D(key[14]), .SP(n68[3]), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key_r[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_r_i14.GSR = "ENABLED";
    LUT4 or_22_i3_2_lut (.A(key_r[6]), .B(key[6]), .Z(key_out_15__N_117[2])) /* synthesis lut_function=(A+(B)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(89[37:60])
    defparam or_22_i3_2_lut.init = 16'heeee;
    FD1S3DX cnt_115_116__i1 (.D(n82[0]), .CK(clk_c), .CD(rst_n_N_6), .Q(\cnt[0] )) /* synthesis syn_use_carry_chain=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(55[12:22])
    defparam cnt_115_116__i1.GSR = "ENABLED";
    LUT4 or_21_i1_2_lut (.A(key_r[0]), .B(key[0]), .Z(key_out_15__N_121[0])) /* synthesis lut_function=(A+(B)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(88[37:60])
    defparam or_21_i1_2_lut.init = 16'heeee;
    FD1S3DX c_state_FSM_i1 (.D(n68[0]), .CK(clk_200hz), .CD(rst_n_N_6), 
            .Q(n68[1]));   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(68[4] 75[11])
    defparam c_state_FSM_i1.GSR = "ENABLED";
    LUT4 i167_2_lut_3_lut (.A(n68[2]), .B(n68[3]), .C(n68[1]), .Z(clk_200hz_N_24_enable_46)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(68[4] 75[11])
    defparam i167_2_lut_3_lut.init = 16'h1010;
    LUT4 or_22_i2_2_lut (.A(key_r[5]), .B(key[5]), .Z(key_out_15__N_117[1])) /* synthesis lut_function=(A+(B)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(89[37:60])
    defparam or_22_i2_2_lut.init = 16'heeee;
    FD1S3DX c_state_FSM_i2 (.D(n68[1]), .CK(clk_200hz), .CD(rst_n_N_6), 
            .Q(n68[2]));   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(68[4] 75[11])
    defparam c_state_FSM_i2.GSR = "ENABLED";
    LUT4 key_out_r_15__I_0_i11_2_lut (.A(key_out_r[10]), .B(key_out[10]), 
         .Z(key_pulse[10])) /* synthesis lut_function=(!((B)+!A)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(105[20:43])
    defparam key_out_r_15__I_0_i11_2_lut.init = 16'h2222;
    LUT4 key_out_r_15__I_0_i9_2_lut (.A(key_out_r[8]), .B(key_out[8]), .Z(key_pulse[8])) /* synthesis lut_function=(!((B)+!A)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(105[20:43])
    defparam key_out_r_15__I_0_i9_2_lut.init = 16'h2222;
    LUT4 i3_2_lut_3_lut (.A(n5), .B(\cnt[13] ), .C(\cnt[12] ), .Z(clk_200hz_N_26)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i3_2_lut_3_lut.init = 16'h8080;
    FD1P3BX key_out_i7 (.D(key_out_15__N_117[3]), .SP(clk_200hz_N_24_enable_46), 
            .CK(clk_200hz_N_24), .PD(rst_n_N_6), .Q(\key_out[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_out_i7.GSR = "ENABLED";
    FD1P3BX key_r_i13 (.D(key[13]), .SP(n68[3]), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key_r[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_r_i13.GSR = "ENABLED";
    FD1P3BX key_r_i12 (.D(key[12]), .SP(n68[3]), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key_r[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_r_i12.GSR = "ENABLED";
    LUT4 key_out_r_15__I_0_i10_2_lut (.A(\key_out_r[9] ), .B(\key_out[9] ), 
         .Z(key_pulse[9])) /* synthesis lut_function=(!((B)+!A)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(105[20:43])
    defparam key_out_r_15__I_0_i10_2_lut.init = 16'h2222;
    FD1S3BX c_state_FSM_i0 (.D(n68[3]), .CK(clk_200hz), .PD(rst_n_N_6), 
            .Q(n68[0]));   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(68[4] 75[11])
    defparam c_state_FSM_i0.GSR = "ENABLED";
    LUT4 or_21_i4_2_lut (.A(key_r[3]), .B(key[3]), .Z(key_out_15__N_121[3])) /* synthesis lut_function=(A+(B)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(88[37:60])
    defparam or_21_i4_2_lut.init = 16'heeee;
    LUT4 key_out_r_15__I_0_i3_2_lut (.A(key_out_r[2]), .B(key_out[2]), .Z(key_pulse[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(105[20:43])
    defparam key_out_r_15__I_0_i3_2_lut.init = 16'h2222;
    LUT4 i169_2_lut_3_lut (.A(n68[2]), .B(n68[3]), .C(n68[1]), .Z(row_3__N_1[1])) /* synthesis lut_function=(A+(B+(C))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(68[4] 75[11])
    defparam i169_2_lut_3_lut.init = 16'hfefe;
    LUT4 or_23_i2_2_lut (.A(key_r[9]), .B(key[9]), .Z(key_out_15__N_113[1])) /* synthesis lut_function=(A+(B)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(90[37:60])
    defparam or_23_i2_2_lut.init = 16'heeee;
    FD1P3BX key_out_i6 (.D(key_out_15__N_117[2]), .SP(clk_200hz_N_24_enable_46), 
            .CK(clk_200hz_N_24), .PD(rst_n_N_6), .Q(\key_out[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_out_i6.GSR = "ENABLED";
    LUT4 key_out_r_15__I_0_i12_2_lut (.A(\key_out_r[11] ), .B(\key_out[11] ), 
         .Z(key_pulse[11])) /* synthesis lut_function=(!((B)+!A)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(105[20:43])
    defparam key_out_r_15__I_0_i12_2_lut.init = 16'h2222;
    FD1P3BX key_r_i11 (.D(key[11]), .SP(clk_200hz_N_24_enable_45), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key_r[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_r_i11.GSR = "ENABLED";
    FD1P3BX key_out_i5 (.D(key_out_15__N_117[1]), .SP(clk_200hz_N_24_enable_46), 
            .CK(clk_200hz_N_24), .PD(rst_n_N_6), .Q(\key_out[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_out_i5.GSR = "ENABLED";
    LUT4 key_out_r_15__I_0_i4_2_lut (.A(key_out_r[3]), .B(key_out[3]), .Z(key_pulse[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(105[20:43])
    defparam key_out_r_15__I_0_i4_2_lut.init = 16'h2222;
    LUT4 i268_2_lut (.A(n68[3]), .B(n68[2]), .Z(row_3__N_1[3])) /* synthesis lut_function=(A+!(B)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(68[4] 75[11])
    defparam i268_2_lut.init = 16'hbbbb;
    LUT4 or_23_i1_2_lut (.A(key_r[8]), .B(key[8]), .Z(key_out_15__N_113[0])) /* synthesis lut_function=(A+(B)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(90[37:60])
    defparam or_23_i1_2_lut.init = 16'heeee;
    LUT4 i1_4_lut (.A(n20), .B(cnt[14]), .C(cnt[11]), .D(cnt[10]), .Z(n5)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i1_4_lut.init = 16'hc8c0;
    LUT4 i149_4_lut (.A(cnt[7]), .B(cnt[9]), .C(cnt[8]), .D(n4), .Z(n20)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;
    defparam i149_4_lut.init = 16'hfcec;
    LUT4 or_22_i1_2_lut (.A(key_r[4]), .B(key[4]), .Z(key_out_15__N_117[0])) /* synthesis lut_function=(A+(B)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(89[37:60])
    defparam or_22_i1_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_2 (.A(cnt[6]), .B(n1047), .C(cnt[5]), .D(cnt[4]), 
         .Z(n4)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_2.init = 16'hfaea;
    LUT4 i366_1_lut_2_lut (.A(n68[3]), .B(n68[2]), .Z(clk_200hz_N_24_enable_45)) /* synthesis lut_function=(!(A+!(B))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(68[4] 75[11])
    defparam i366_1_lut_2_lut.init = 16'h4444;
    LUT4 key_out_r_15__I_0_i15_2_lut (.A(key_out_r[14]), .B(key_out[14]), 
         .Z(key_pulse[14])) /* synthesis lut_function=(!((B)+!A)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(105[20:43])
    defparam key_out_r_15__I_0_i15_2_lut.init = 16'h2222;
    LUT4 key_out_r_15__I_0_i1_2_lut (.A(\key_out_r[0] ), .B(\key_out[0] ), 
         .Z(key_pulse[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(105[20:43])
    defparam key_out_r_15__I_0_i1_2_lut.init = 16'h2222;
    FD1P3BX key_out_i4 (.D(key_out_15__N_117[0]), .SP(clk_200hz_N_24_enable_46), 
            .CK(clk_200hz_N_24), .PD(rst_n_N_6), .Q(\key_out[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_out_i4.GSR = "ENABLED";
    FD1P3BX key_r_i10 (.D(key[10]), .SP(clk_200hz_N_24_enable_45), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key_r[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_r_i10.GSR = "ENABLED";
    FD1P3BX key_r_i9 (.D(key[9]), .SP(clk_200hz_N_24_enable_45), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key_r[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_r_i9.GSR = "ENABLED";
    LUT4 key_out_r_15__I_0_i2_2_lut (.A(\key_out_r[1] ), .B(\key_out[1] ), 
         .Z(key_pulse[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(105[20:43])
    defparam key_out_r_15__I_0_i2_2_lut.init = 16'h2222;
    FD1P3BX key_r_i8 (.D(key[8]), .SP(clk_200hz_N_24_enable_45), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key_r[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_r_i8.GSR = "ENABLED";
    LUT4 key_out_r_15__I_0_i5_2_lut (.A(\key_out_r[4] ), .B(\key_out[4] ), 
         .Z(key_pulse[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(105[20:43])
    defparam key_out_r_15__I_0_i5_2_lut.init = 16'h2222;
    LUT4 i3_4_lut (.A(\cnt[0] ), .B(cnt[3]), .C(cnt[2]), .D(cnt[1]), 
         .Z(n1047)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 key_out_r_15__I_0_i16_2_lut (.A(\key_out_r[15] ), .B(\key_out[15] ), 
         .Z(key_pulse[15])) /* synthesis lut_function=(!((B)+!A)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(105[20:43])
    defparam key_out_r_15__I_0_i16_2_lut.init = 16'h2222;
    LUT4 i2_2_lut (.A(\cnt[13] ), .B(\cnt[12] ), .Z(n6)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 key_out_r_15__I_0_i6_2_lut (.A(\key_out_r[5] ), .B(\key_out[5] ), 
         .Z(key_pulse[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(105[20:43])
    defparam key_out_r_15__I_0_i6_2_lut.init = 16'h2222;
    LUT4 i445_2_lut_3_lut (.A(n68[2]), .B(n68[3]), .C(n68[1]), .Z(row_3__N_1[2])) /* synthesis lut_function=(A+(B+!(C))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(68[4] 75[11])
    defparam i445_2_lut_3_lut.init = 16'hefef;
    LUT4 or_21_i3_2_lut (.A(key_r[2]), .B(key[2]), .Z(key_out_15__N_121[2])) /* synthesis lut_function=(A+(B)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(88[37:60])
    defparam or_21_i3_2_lut.init = 16'heeee;
    FD1P3BX key_r_i7 (.D(key[7]), .SP(clk_200hz_N_24_enable_46), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key_r[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_r_i7.GSR = "ENABLED";
    LUT4 i77_1_lut (.A(n68[3]), .Z(row_3__N_1[0])) /* synthesis lut_function=(!(A)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(68[4] 75[11])
    defparam i77_1_lut.init = 16'h5555;
    LUT4 clk_200hz_I_0_47_2_lut_3_lut_4_lut (.A(clk_200hz), .B(n5), .C(\cnt[13] ), 
         .D(\cnt[12] ), .Z(clk_200hz_N_25)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B (C (D))))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(54[13] 57[7])
    defparam clk_200hz_I_0_47_2_lut_3_lut_4_lut.init = 16'h6aaa;
    LUT4 or_21_i2_2_lut (.A(key_r[1]), .B(key[1]), .Z(key_out_15__N_121[1])) /* synthesis lut_function=(A+(B)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(88[37:60])
    defparam or_21_i2_2_lut.init = 16'heeee;
    FD1P3BX key_out_i3 (.D(key_out_15__N_121[3]), .SP(clk_200hz_N_24_enable_48), 
            .CK(clk_200hz_N_24), .PD(rst_n_N_6), .Q(key_out[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_out_i3.GSR = "ENABLED";
    CCU2D cnt_115_116_add_4_15 (.A0(\cnt[13] ), .B0(clk_200hz_N_26), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[14]), .B1(clk_200hz_N_26), .C1(GND_net), 
          .D1(GND_net), .CIN(n1040), .S0(n82[13]), .S1(n82[14]));   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(55[12:22])
    defparam cnt_115_116_add_4_15.INIT0 = 16'hd222;
    defparam cnt_115_116_add_4_15.INIT1 = 16'hd222;
    defparam cnt_115_116_add_4_15.INJECT1_0 = "NO";
    defparam cnt_115_116_add_4_15.INJECT1_1 = "NO";
    CCU2D cnt_115_116_add_4_13 (.A0(cnt[11]), .B0(clk_200hz_N_26), .C0(GND_net), 
          .D0(GND_net), .A1(\cnt[12] ), .B1(clk_200hz_N_26), .C1(GND_net), 
          .D1(GND_net), .CIN(n1039), .COUT(n1040), .S0(n82[11]), .S1(n82[12]));   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(55[12:22])
    defparam cnt_115_116_add_4_13.INIT0 = 16'hd222;
    defparam cnt_115_116_add_4_13.INIT1 = 16'hd222;
    defparam cnt_115_116_add_4_13.INJECT1_0 = "NO";
    defparam cnt_115_116_add_4_13.INJECT1_1 = "NO";
    CCU2D cnt_115_116_add_4_11 (.A0(cnt[9]), .B0(clk_200hz_N_26), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[10]), .B1(clk_200hz_N_26), .C1(GND_net), 
          .D1(GND_net), .CIN(n1038), .COUT(n1039), .S0(n82[9]), .S1(n82[10]));   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(55[12:22])
    defparam cnt_115_116_add_4_11.INIT0 = 16'hd222;
    defparam cnt_115_116_add_4_11.INIT1 = 16'hd222;
    defparam cnt_115_116_add_4_11.INJECT1_0 = "NO";
    defparam cnt_115_116_add_4_11.INJECT1_1 = "NO";
    CCU2D cnt_115_116_add_4_9 (.A0(cnt[7]), .B0(clk_200hz_N_26), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[8]), .B1(clk_200hz_N_26), .C1(GND_net), 
          .D1(GND_net), .CIN(n1037), .COUT(n1038), .S0(n82[7]), .S1(n82[8]));   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(55[12:22])
    defparam cnt_115_116_add_4_9.INIT0 = 16'hd222;
    defparam cnt_115_116_add_4_9.INIT1 = 16'hd222;
    defparam cnt_115_116_add_4_9.INJECT1_0 = "NO";
    defparam cnt_115_116_add_4_9.INJECT1_1 = "NO";
    CCU2D cnt_115_116_add_4_7 (.A0(cnt[5]), .B0(clk_200hz_N_26), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[6]), .B1(clk_200hz_N_26), .C1(GND_net), 
          .D1(GND_net), .CIN(n1036), .COUT(n1037), .S0(n82[5]), .S1(n82[6]));   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(55[12:22])
    defparam cnt_115_116_add_4_7.INIT0 = 16'hd222;
    defparam cnt_115_116_add_4_7.INIT1 = 16'hd222;
    defparam cnt_115_116_add_4_7.INJECT1_0 = "NO";
    defparam cnt_115_116_add_4_7.INJECT1_1 = "NO";
    CCU2D cnt_115_116_add_4_5 (.A0(cnt[3]), .B0(clk_200hz_N_26), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[4]), .B1(clk_200hz_N_26), .C1(GND_net), 
          .D1(GND_net), .CIN(n1035), .COUT(n1036), .S0(n82[3]), .S1(n82[4]));   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(55[12:22])
    defparam cnt_115_116_add_4_5.INIT0 = 16'hd222;
    defparam cnt_115_116_add_4_5.INIT1 = 16'hd222;
    defparam cnt_115_116_add_4_5.INJECT1_0 = "NO";
    defparam cnt_115_116_add_4_5.INJECT1_1 = "NO";
    CCU2D cnt_115_116_add_4_3 (.A0(cnt[1]), .B0(clk_200hz_N_26), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[2]), .B1(clk_200hz_N_26), .C1(GND_net), 
          .D1(GND_net), .CIN(n1034), .COUT(n1035), .S0(n82[1]), .S1(n82[2]));   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(55[12:22])
    defparam cnt_115_116_add_4_3.INIT0 = 16'hd222;
    defparam cnt_115_116_add_4_3.INIT1 = 16'hd222;
    defparam cnt_115_116_add_4_3.INJECT1_0 = "NO";
    defparam cnt_115_116_add_4_3.INJECT1_1 = "NO";
    FD1P3BX key_out_i2 (.D(key_out_15__N_121[2]), .SP(clk_200hz_N_24_enable_48), 
            .CK(clk_200hz_N_24), .PD(rst_n_N_6), .Q(key_out[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_out_i2.GSR = "ENABLED";
    FD1P3BX key_r_i6 (.D(key[6]), .SP(clk_200hz_N_24_enable_46), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key_r[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_r_i6.GSR = "ENABLED";
    FD1P3BX key_r_i5 (.D(key[5]), .SP(clk_200hz_N_24_enable_46), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key_r[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_r_i5.GSR = "ENABLED";
    LUT4 or_24_i4_2_lut (.A(key_r[15]), .B(key[15]), .Z(key_out_15__N_109[3])) /* synthesis lut_function=(A+(B)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(91[37:60])
    defparam or_24_i4_2_lut.init = 16'heeee;
    OFS1P3BX row_i3 (.D(row_3__N_1[2]), .SP(VCC_net), .SCLK(clk_200hz), 
            .PD(rst_n_N_6), .Q(row_c_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(67[12] 76[6])
    defparam row_i3.GSR = "ENABLED";
    OFS1P3BX row_i2 (.D(row_3__N_1[1]), .SP(VCC_net), .SCLK(clk_200hz), 
            .PD(rst_n_N_6), .Q(row_c_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(67[12] 76[6])
    defparam row_i2.GSR = "ENABLED";
    FD1S3DX cnt_115_116__i15 (.D(n82[14]), .CK(clk_c), .CD(rst_n_N_6), 
            .Q(cnt[14])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(55[12:22])
    defparam cnt_115_116__i15.GSR = "ENABLED";
    OFS1P3DX row_i1 (.D(row_3__N_1[0]), .SP(VCC_net), .SCLK(clk_200hz), 
            .CD(rst_n_N_6), .Q(row_c_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(67[12] 76[6])
    defparam row_i1.GSR = "ENABLED";
    CCU2D cnt_115_116_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n5), .B1(n6), .C1(n1032), .D1(GND_net), 
          .COUT(n1034), .S1(n82[0]));   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(55[12:22])
    defparam cnt_115_116_add_4_1.INIT0 = 16'hF000;
    defparam cnt_115_116_add_4_1.INIT1 = 16'h8787;
    defparam cnt_115_116_add_4_1.INJECT1_0 = "NO";
    defparam cnt_115_116_add_4_1.INJECT1_1 = "NO";
    FD1S3DX cnt_115_116__i14 (.D(n82[13]), .CK(clk_c), .CD(rst_n_N_6), 
            .Q(\cnt[13] )) /* synthesis syn_use_carry_chain=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(55[12:22])
    defparam cnt_115_116__i14.GSR = "ENABLED";
    FD1S3DX cnt_115_116__i13 (.D(n82[12]), .CK(clk_c), .CD(rst_n_N_6), 
            .Q(\cnt[12] )) /* synthesis syn_use_carry_chain=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(55[12:22])
    defparam cnt_115_116__i13.GSR = "ENABLED";
    FD1S3DX cnt_115_116__i12 (.D(n82[11]), .CK(clk_c), .CD(rst_n_N_6), 
            .Q(cnt[11])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(55[12:22])
    defparam cnt_115_116__i12.GSR = "ENABLED";
    FD1S3DX cnt_115_116__i11 (.D(n82[10]), .CK(clk_c), .CD(rst_n_N_6), 
            .Q(cnt[10])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(55[12:22])
    defparam cnt_115_116__i11.GSR = "ENABLED";
    FD1S3DX cnt_115_116__i10 (.D(n82[9]), .CK(clk_c), .CD(rst_n_N_6), 
            .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(55[12:22])
    defparam cnt_115_116__i10.GSR = "ENABLED";
    FD1S3DX cnt_115_116__i9 (.D(n82[8]), .CK(clk_c), .CD(rst_n_N_6), .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(55[12:22])
    defparam cnt_115_116__i9.GSR = "ENABLED";
    FD1S3DX cnt_115_116__i8 (.D(n82[7]), .CK(clk_c), .CD(rst_n_N_6), .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(55[12:22])
    defparam cnt_115_116__i8.GSR = "ENABLED";
    FD1S3DX cnt_115_116__i7 (.D(n82[6]), .CK(clk_c), .CD(rst_n_N_6), .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(55[12:22])
    defparam cnt_115_116__i7.GSR = "ENABLED";
    FD1S3BX key_out_r_i15 (.D(\key_out[15] ), .CK(clk_c), .PD(rst_n_N_6), 
            .Q(\key_out_r[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(101[9:30])
    defparam key_out_r_i15.GSR = "ENABLED";
    FD1P3BX key_r_i4 (.D(key[4]), .SP(clk_200hz_N_24_enable_46), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key_r[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_r_i4.GSR = "ENABLED";
    FD1P3BX key_r_i3 (.D(key[3]), .SP(clk_200hz_N_24_enable_48), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key_r[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_r_i3.GSR = "ENABLED";
    FD1S3BX key_out_r_i14 (.D(key_out[14]), .CK(clk_c), .PD(rst_n_N_6), 
            .Q(key_out_r[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(101[9:30])
    defparam key_out_r_i14.GSR = "ENABLED";
    FD1S3BX key_out_r_i13 (.D(\key_out[13] ), .CK(clk_c), .PD(rst_n_N_6), 
            .Q(\key_out_r[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(101[9:30])
    defparam key_out_r_i13.GSR = "ENABLED";
    FD1S3BX key_out_r_i12 (.D(key_out[12]), .CK(clk_c), .PD(rst_n_N_6), 
            .Q(key_out_r[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(101[9:30])
    defparam key_out_r_i12.GSR = "ENABLED";
    FD1S3BX key_out_r_i11 (.D(\key_out[11] ), .CK(clk_c), .PD(rst_n_N_6), 
            .Q(\key_out_r[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(101[9:30])
    defparam key_out_r_i11.GSR = "ENABLED";
    FD1S3DX cnt_115_116__i6 (.D(n82[5]), .CK(clk_c), .CD(rst_n_N_6), .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(55[12:22])
    defparam cnt_115_116__i6.GSR = "ENABLED";
    FD1S3DX cnt_115_116__i5 (.D(n82[4]), .CK(clk_c), .CD(rst_n_N_6), .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(55[12:22])
    defparam cnt_115_116__i5.GSR = "ENABLED";
    FD1S3DX cnt_115_116__i4 (.D(n82[3]), .CK(clk_c), .CD(rst_n_N_6), .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(55[12:22])
    defparam cnt_115_116__i4.GSR = "ENABLED";
    FD1S3BX key_out_r_i10 (.D(key_out[10]), .CK(clk_c), .PD(rst_n_N_6), 
            .Q(key_out_r[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(101[9:30])
    defparam key_out_r_i10.GSR = "ENABLED";
    FD1S3BX key_out_r_i9 (.D(\key_out[9] ), .CK(clk_c), .PD(rst_n_N_6), 
            .Q(\key_out_r[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(101[9:30])
    defparam key_out_r_i9.GSR = "ENABLED";
    FD1S3BX key_out_r_i8 (.D(key_out[8]), .CK(clk_c), .PD(rst_n_N_6), 
            .Q(key_out_r[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(101[9:30])
    defparam key_out_r_i8.GSR = "ENABLED";
    FD1S3BX key_out_r_i7 (.D(\key_out[7] ), .CK(clk_c), .PD(rst_n_N_6), 
            .Q(\key_out_r[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(101[9:30])
    defparam key_out_r_i7.GSR = "ENABLED";
    FD1S3BX key_out_r_i6 (.D(\key_out[6] ), .CK(clk_c), .PD(rst_n_N_6), 
            .Q(\key_out_r[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(101[9:30])
    defparam key_out_r_i6.GSR = "ENABLED";
    FD1S3BX key_out_r_i5 (.D(\key_out[5] ), .CK(clk_c), .PD(rst_n_N_6), 
            .Q(\key_out_r[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(101[9:30])
    defparam key_out_r_i5.GSR = "ENABLED";
    FD1S3BX key_out_r_i4 (.D(\key_out[4] ), .CK(clk_c), .PD(rst_n_N_6), 
            .Q(\key_out_r[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(101[9:30])
    defparam key_out_r_i4.GSR = "ENABLED";
    FD1S3BX key_out_r_i3 (.D(key_out[3]), .CK(clk_c), .PD(rst_n_N_6), 
            .Q(key_out_r[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(101[9:30])
    defparam key_out_r_i3.GSR = "ENABLED";
    FD1S3DX cnt_115_116__i3 (.D(n82[2]), .CK(clk_c), .CD(rst_n_N_6), .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(55[12:22])
    defparam cnt_115_116__i3.GSR = "ENABLED";
    FD1S3DX cnt_115_116__i2 (.D(n82[1]), .CK(clk_c), .CD(rst_n_N_6), .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(55[12:22])
    defparam cnt_115_116__i2.GSR = "ENABLED";
    FD1P3BX key_out_i1 (.D(key_out_15__N_121[1]), .SP(clk_200hz_N_24_enable_48), 
            .CK(clk_200hz_N_24), .PD(rst_n_N_6), .Q(\key_out[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_out_i1.GSR = "ENABLED";
    LUT4 i365_1_lut_3_lut (.A(n68[2]), .B(n68[3]), .C(n68[1]), .Z(clk_200hz_N_24_enable_48)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(68[4] 75[11])
    defparam i365_1_lut_3_lut.init = 16'h0101;
    LUT4 or_24_i3_2_lut (.A(key_r[14]), .B(key[14]), .Z(key_out_15__N_109[2])) /* synthesis lut_function=(A+(B)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(91[37:60])
    defparam or_24_i3_2_lut.init = 16'heeee;
    LUT4 key_out_r_15__I_0_i7_2_lut (.A(\key_out_r[6] ), .B(\key_out[6] ), 
         .Z(key_pulse[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(105[20:43])
    defparam key_out_r_15__I_0_i7_2_lut.init = 16'h2222;
    FD1S3DX c_state_FSM_i3 (.D(n68[2]), .CK(clk_200hz), .CD(rst_n_N_6), 
            .Q(n68[3]));   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(68[4] 75[11])
    defparam c_state_FSM_i3.GSR = "ENABLED";
    FD1P3BX key_r_i2 (.D(key[2]), .SP(clk_200hz_N_24_enable_48), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key_r[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_r_i2.GSR = "ENABLED";
    FD1S3BX key_out_r_i2 (.D(key_out[2]), .CK(clk_c), .PD(rst_n_N_6), 
            .Q(key_out_r[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(101[9:30])
    defparam key_out_r_i2.GSR = "ENABLED";
    FD1S3BX key_out_r_i1 (.D(\key_out[1] ), .CK(clk_c), .PD(rst_n_N_6), 
            .Q(\key_out_r[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(101[9:30])
    defparam key_out_r_i1.GSR = "ENABLED";
    FD1P3BX key_i15 (.D(col_c_3), .SP(n68[3]), .CK(clk_200hz_N_24), .PD(rst_n_N_6), 
            .Q(key[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_i15.GSR = "ENABLED";
    FD1P3BX key_r_i1 (.D(key[1]), .SP(clk_200hz_N_24_enable_48), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key_r[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_r_i1.GSR = "ENABLED";
    FD1P3BX key_i14 (.D(col_c_2), .SP(n68[3]), .CK(clk_200hz_N_24), .PD(rst_n_N_6), 
            .Q(key[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_i14.GSR = "ENABLED";
    FD1P3BX key_out_i15 (.D(key_out_15__N_109[3]), .SP(n68[3]), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(\key_out[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_out_i15.GSR = "ENABLED";
    OFS1P3BX row_i4 (.D(row_3__N_1[3]), .SP(VCC_net), .SCLK(clk_200hz), 
            .PD(rst_n_N_6), .Q(row_c_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(67[12] 76[6])
    defparam row_i4.GSR = "ENABLED";
    FD1P3BX key_i13 (.D(col_c_1), .SP(n68[3]), .CK(clk_200hz_N_24), .PD(rst_n_N_6), 
            .Q(key[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_i13.GSR = "ENABLED";
    FD1P3BX key_i12 (.D(col_c_0), .SP(n68[3]), .CK(clk_200hz_N_24), .PD(rst_n_N_6), 
            .Q(key[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_i12.GSR = "ENABLED";
    FD1P3BX key_out_i14 (.D(key_out_15__N_109[2]), .SP(n68[3]), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key_out[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_out_i14.GSR = "ENABLED";
    FD1P3BX key_i11 (.D(col_c_3), .SP(clk_200hz_N_24_enable_45), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_i11.GSR = "ENABLED";
    LUT4 or_24_i2_2_lut (.A(key_r[13]), .B(key[13]), .Z(key_out_15__N_109[1])) /* synthesis lut_function=(A+(B)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(91[37:60])
    defparam or_24_i2_2_lut.init = 16'heeee;
    FD1P3BX key_out_i13 (.D(key_out_15__N_109[1]), .SP(n68[3]), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(\key_out[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_out_i13.GSR = "ENABLED";
    LUT4 or_24_i1_2_lut (.A(key_r[12]), .B(key[12]), .Z(key_out_15__N_109[0])) /* synthesis lut_function=(A+(B)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(91[37:60])
    defparam or_24_i1_2_lut.init = 16'heeee;
    FD1P3BX key_i10 (.D(col_c_2), .SP(clk_200hz_N_24_enable_45), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_i10.GSR = "ENABLED";
    FD1P3BX key_i9 (.D(col_c_1), .SP(clk_200hz_N_24_enable_45), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_i9.GSR = "ENABLED";
    LUT4 key_out_r_15__I_0_i8_2_lut (.A(\key_out_r[7] ), .B(\key_out[7] ), 
         .Z(key_pulse[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(105[20:43])
    defparam key_out_r_15__I_0_i8_2_lut.init = 16'h2222;
    FD1P3BX key_out_i12 (.D(key_out_15__N_109[0]), .SP(n68[3]), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key_out[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_out_i12.GSR = "ENABLED";
    FD1P3BX key_out_i11 (.D(key_out_15__N_113[3]), .SP(clk_200hz_N_24_enable_45), 
            .CK(clk_200hz_N_24), .PD(rst_n_N_6), .Q(\key_out[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_out_i11.GSR = "ENABLED";
    FD1P3BX key_i8 (.D(col_c_0), .SP(clk_200hz_N_24_enable_45), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_i8.GSR = "ENABLED";
    FD1P3BX key_i7 (.D(col_c_3), .SP(clk_200hz_N_24_enable_46), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_i7.GSR = "ENABLED";
    FD1P3BX key_i6 (.D(col_c_2), .SP(clk_200hz_N_24_enable_46), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_i6.GSR = "ENABLED";
    FD1P3BX key_i5 (.D(col_c_1), .SP(clk_200hz_N_24_enable_46), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_i5.GSR = "ENABLED";
    FD1P3BX key_out_i10 (.D(key_out_15__N_113[2]), .SP(clk_200hz_N_24_enable_45), 
            .CK(clk_200hz_N_24), .PD(rst_n_N_6), .Q(key_out[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_out_i10.GSR = "ENABLED";
    FD1P3BX key_i4 (.D(col_c_0), .SP(clk_200hz_N_24_enable_46), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_i4.GSR = "ENABLED";
    FD1P3BX key_i3 (.D(col_c_3), .SP(clk_200hz_N_24_enable_48), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_i3.GSR = "ENABLED";
    LUT4 or_23_i4_2_lut (.A(key_r[11]), .B(key[11]), .Z(key_out_15__N_113[3])) /* synthesis lut_function=(A+(B)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(90[37:60])
    defparam or_23_i4_2_lut.init = 16'heeee;
    LUT4 or_23_i3_2_lut (.A(key_r[10]), .B(key[10]), .Z(key_out_15__N_113[2])) /* synthesis lut_function=(A+(B)) */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(90[37:60])
    defparam or_23_i3_2_lut.init = 16'heeee;
    FD1P3BX key_i2 (.D(col_c_2), .SP(clk_200hz_N_24_enable_48), .CK(clk_200hz_N_24), 
            .PD(rst_n_N_6), .Q(key[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=31, LSE_RLINE=39 */ ;   // f:/fpga_project/baseboard/lab1_type_system/array_keyboard.v(84[12] 94[6])
    defparam key_i2.GSR = "ENABLED";
    
endmodule
