`timescale 1ns / 100ps
module step_rom (Address, Q);

    input wire [6:0] Address;
    output reg [127:0] Q;
	 
	always @ (*)
		case(Address)
			8'd0  : Q = 128'h00000000000000000000000000000000;
			8'd1  : Q = 128'h00000000000000000000000000000000;
			8'd2  : Q = 128'h00000000000000000000000000000000;
			8'd3  : Q = 128'h000000000000001C0000000000000000;
			8'd4  : Q = 128'h00000000000001FFC000000000000000;
			8'd5  : Q = 128'h00000000000003FFE000000000000000;
			8'd6  : Q = 128'h00000000000007FFF800000000000000;
			8'd7  : Q = 128'h0000000000001FFFFC00000000000000;
			8'd8  : Q = 128'h0000000000003FFFFF00000000000000;
			8'd9  : Q = 128'h0000000000007FFFFF80000000000000;
			8'd10 : Q = 128'h000000000000FFFFFF80000000000000;
			8'd11 : Q = 128'h000000000000FFFFFFC0000000000000;
			8'd12 : Q = 128'h000000000001FFFFFFC0000000000000;
			8'd13 : Q = 128'h000000000001FFFFFFE0000000000000;
			8'd14 : Q = 128'h000000000003FFFFFFE0000000000000;
			8'd15 : Q = 128'h000000000003FFFFFFE0000000000000;
			8'd16 : Q = 128'h000000000007FFC1FFF0000000000000;
			8'd17 : Q = 128'h000000000007FF807FF0000000000000;
			8'd18 : Q = 128'h000000000007FF007FF0000000000000;
			8'd19 : Q = 128'h000000000007FF007FF0000000000000;
			8'd20 : Q = 128'h000000000007FF007FF0000000000000;
			8'd21 : Q = 128'h000000000007FF007FF0000000000000;
			8'd22 : Q = 128'h000000000007FF80FFF0000000000000;
			8'd23 : Q = 128'h000000000007FF81FFF0000000000000;
			8'd24 : Q = 128'h000000000007FFC3FFE0000000000000;
			8'd25 : Q = 128'h000000000003FFE7FFE0000000000000;
			8'd26 : Q = 128'h000000000001FFE7FFE0000000000000;
			8'd27 : Q = 128'h000000000001FFE7FFC00000007FC000;
			8'd28 : Q = 128'h000000000000FFE7FFC0000001FFF000;
			8'd29 : Q = 128'h000000000000FFE7FF80000007FFFC00;
			8'd30 : Q = 128'h000FF80000007FE7FF0000001FFFFF00;
			8'd31 : Q = 128'h003FFE0000007FE7FF0000003FFFFF80;
			8'd32 : Q = 128'h00FFFE0000007FE7FE0000003FFFFF80;
			8'd33 : Q = 128'h01FFFF0000003FE7FE0000007FFFFFC0;
			8'd34 : Q = 128'h03FFFF8000003FE7FC0000007FFFFFC0;
			8'd35 : Q = 128'h07FFFFE000001FCFFC000000FFFFFFE0;
			8'd36 : Q = 128'h07FFFFF000001FCFFC000000FFFFFFE0;
			8'd37 : Q = 128'h0FFFFFF000001FCFF8000000FFF9FFE0;
			8'd38 : Q = 128'h0FFF7FF800000FCFF8000001FFE07FF0;
			8'd39 : Q = 128'h0FFC1FF800000FCFF0000001FFE07FF0;
			8'd40 : Q = 128'h1FF80FF800000FCFF0000001FFC03FF0;
			8'd41 : Q = 128'h1FF80FF800000FCFF0000001FFC03FF0;
			8'd42 : Q = 128'h1FF00FF800000FCFF0000001FFC03FF0;
			8'd43 : Q = 128'h1FF00FF800000FCFE0000001FFC03FF0;
			8'd44 : Q = 128'h1FF80FFC00000FCFE0000001FFE07FF0;
			8'd45 : Q = 128'h0FF81FF8000007CFE0000003FFC0FFE0;
			8'd46 : Q = 128'h0FFC1FF8000007CFE0000003FF87FFE0;
			8'd47 : Q = 128'h0FFF8FF8000007CFC0000003FF8FFFE0;
			8'd48 : Q = 128'h0FFF8FF80000079FC0000003FF1FFFC0;
			8'd49 : Q = 128'h07FFCFF80000079FC0000007FF3FFFC0;
			8'd50 : Q = 128'h07FFCFF80000079FC0000007FE3FFF80;
			8'd51 : Q = 128'h03FFC7F80000079FC0000007FC7FFF80;
			8'd52 : Q = 128'h03FFE7F80000079FC0000007F8FFFF00;
			8'd53 : Q = 128'h01FFE3FC0000079F8000000FF0FFFC00;
			8'd54 : Q = 128'h007FF3FC0000079F8000000FE1FFF800;
			8'd55 : Q = 128'h001FF3FC0000079F8000001FC3FFF000;
			8'd56 : Q = 128'h0007F9FC0000079F8000001F8FFFC000;
			8'd57 : Q = 128'h0003F9FC0000071F8000003F9FFF8000;
			8'd58 : Q = 128'h0001F8FC00000F3F8000003F1FFF0000;
			8'd59 : Q = 128'h0000FCFC00000F3F8000003F3FFE0000;
			8'd60 : Q = 128'h00007CFC00000F3F8000007E3FFC0000;
			8'd61 : Q = 128'h00003E7C00000F3F8000007C7FF80000;
			8'd62 : Q = 128'h00001E7E00000F3F800000F8FFE00000;
			8'd63 : Q = 128'h00001F3E00000F3F800001F1FFC00000;
			8'd64 : Q = 128'h00000F1E00001F3FC00001F3FF800000;
			8'd65 : Q = 128'h0000078F00001F3FC00003E3FE000000;
			8'd66 : Q = 128'h0000078700001E3FE00007C7FC000000;
			8'd67 : Q = 128'h000003C780003E3FF0000F8FF0000000;
			8'd68 : Q = 128'h000003C780003E3FF0001F9FE0000000;
			8'd69 : Q = 128'h000003E3C0007E3FF8001F1FE0000000;
			8'd70 : Q = 128'h000001F3C000FE3FFC007F3FC0000000;
			8'd71 : Q = 128'h000001F1E001FE3FFE01FE7F80000000;
			8'd72 : Q = 128'h000000F9FC0FFC1FFFFFFC7F00000000;
			8'd73 : Q = 128'h000000FCFFFFFC9FFFFFF8FE00000000;
			8'd74 : Q = 128'h0000007C7FFFF88FFFFFF1FC00000000;
			8'd75 : Q = 128'h0000007E3FFFF1CFFFFFC3F800000000;
			8'd76 : Q = 128'h0000003F1FFFF3C7FFFF07F000000000;
			8'd77 : Q = 128'h0000003F8FFFC3E3FFFE0FE000000000;
			8'd78 : Q = 128'h0000003F87FF87F1FFFC1FE000000000;
			8'd79 : Q = 128'h0000001FC1FE0FF07FF87FC000000000;
			8'd80 : Q = 128'h0000000FF0001FFC0FC0FFC000000000;
			8'd81 : Q = 128'h00000007FC00FFFE0003FF8000000000;
			8'd82 : Q = 128'h00000007FFFFFFFFE01FFF0000000000;
			8'd83 : Q = 128'h00000007FFFFFFFFFFFFFF0000000000;
			8'd84 : Q = 128'h00000003FFFFFFFFFFFFFE0000000000;
			8'd85 : Q = 128'h00000003FFFFFFFFFFFFFE0000000000;
			8'd86 : Q = 128'h00000001FFFFFFFFFFFFFC0000000000;
			8'd87 : Q = 128'h00000001FFFFFFFFFFFFFC0000000000;
			8'd88 : Q = 128'h00000001FFFFFFFFFFFFFC0000000000;
			8'd89 : Q = 128'h00000000FFFFFFFFFFFFF80000000000;
			8'd90 : Q = 128'h00000000FFFFFFFFFFFFF80000000000;
			8'd91 : Q = 128'h00000000FFFFFFFFFFFFF00000000000;
			8'd92 : Q = 128'h000000007FFFFFFFFFFFF00000000000;
			8'd93 : Q = 128'h000000007FFFFFFFFFFFE00000000000;
			8'd94 : Q = 128'h000000007FFFFFFFFFFFE00000000000;
			8'd95 : Q = 128'h000000007FFFFFFFFFFFE00000000000;
			8'd96 : Q = 128'h000000003FFFFFFFFFFFC00000000000;
			8'd97 : Q = 128'h000000003FFFFFFFFFFFC00000000000;
			8'd98 : Q = 128'h000000003FFFFFFFFFFF800000000000;
			8'd99 : Q = 128'h000000001FFFFFFFFFFF800000000000;
			8'd100: Q = 128'h000000001FFFFFFFFFFF000000000000;
			8'd101: Q = 128'h000000001FFFFFFFFFFF000000000000;
			8'd102: Q = 128'h000000000FFFFFFFFFFE000000000000;
			8'd103: Q = 128'h000000000FFFFFFFFFFE000000000000;
			8'd104: Q = 128'h000000000FFFFFFFFFFE000000000000;
			8'd105: Q = 128'h000000000FFFFFFFFFFE000000000000;
			8'd106: Q = 128'h0000000007FFFFFFFFFC000000000000;
			8'd107: Q = 128'h0000000007FFFFFFFFFC000000000000;
			8'd108: Q = 128'h0000000007FFFFFFFFFC000000000000;
			8'd109: Q = 128'h0000000003FFFFFFFFF8000000000000;
			8'd110: Q = 128'h0000000003FFFFFFFFF8000000000000;
			8'd111: Q = 128'h0000000001FFFFFFFFF0000000000000;
			8'd112: Q = 128'h0000000000FFFFFFFFE0000000000000;
			8'd113: Q = 128'h0000000000FFFFFFFFE0000000000000;
			8'd114: Q = 128'h0000000000FFFFFFFFC0000000000000;
			8'd115: Q = 128'h00000000007FFFFFFFC0000000000000;
			8'd116: Q = 128'h00000000003FFFFFFF80000000000000;
			8'd117: Q = 128'h00000000001FFFFFFF00000000000000;
			8'd118: Q = 128'h00000000000FFFFFFE00000000000000;
			8'd119: Q = 128'h000000000001FFFFF800000000000000;
			8'd120: Q = 128'h0000000000007FFFE000000000000000;
			8'd121: Q = 128'h0000000000001FFF8000000000000000;
			8'd122: Q = 128'h00000000000003F80000000000000000;
			8'd123: Q = 128'h00000000000000000000000000000000;
			8'd124: Q = 128'h00000000000000000000000000000000;
			8'd125: Q = 128'h00000000000000000000000000000000;
			8'd126: Q = 128'h00000000000000000000000000000000;
			8'd127: Q = 128'h00000000000000000000000000000000;
			default:Q = 128'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
		endcase
		
endmodule
