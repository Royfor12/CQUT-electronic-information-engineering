 // --------------------------------------------------------------------
// >>>>>>>>>>>>>>>>>>>>>>>>> COPYRIGHT NOTICE <<<<<<<<<<<<<<<<<<<<<<<<<
// --------------------------------------------------------------------
// Module: Calculate
// 
// Author: Step
// 
// Description: Calculate
// 
// Web: www.stepfpga.com
// 
// --------------------------------------------------------------------
// Code Revision History :
// --------------------------------------------------------------------
// Version: |Mod. Date:   |Changes Made:
// V1.0     |2016/04/20   |Initial ver
// --------------------------------------------------------------------
module Calculate
(
input				rst_n,		//��λ�ź�
input		[15:0]	T_code,		//�¶���ֵ
input		[15:0]	H_code,		//ʪ����ֵ

output		[15:0]	T_data,		//�¶�BCD��
output		[15:0]	H_data,		//ʪ��BCD��
output		[7:0]	dat_en,		//������ʾʹ��
output		[7:0]	dot_en		//С������ʾʹ��
);

/////////////////////////////////////�¶�����/////////////////////////////////////////

// �¶� T = -46.85 + 175.72 * T_code / 2^16 = (-4685 + 17572 * T_code / 2^16) / 100
wire [31:0] a = T_code * 16'd17572;
wire [31:0] b = a >> 16; //����2^16ȡ��
wire [31:0] c = (b>=32'd4685)? (b - 32'd4685):(32'd4685 - b); //�¶���������ȡ����ֵ
wire [15:0] T_data_bin = c[15:0];

//����BCDת�봦��
//С������BCD�����������2λ����ɳ���100�Ĳ���
//T_data_bcd[19:16]��λ,[15:12]ʮλ,[11:8]��λ,[7:0]����С��λ
wire [19:0] T_data_bcd;
bin_to_bcd u1
(
.rst_n				(rst_n		),	//ϵͳ��λ������Ч
.bin_code			(T_data_bin	),	//��Ҫ����BCDת��Ķ���������
.bcd_code			(T_data_bcd	)	//ת����BCD�����������
);

//Ҫ��ʾ������,����1λС��
//���¶�Ϊ������T_data_bcd[19:16]��λ����������A�滻��ͬʱ�������A���ֿ���ʾ����
assign T_data = (b>=32'd4685)? T_data_bcd[19:4]:{4'ha,T_data_bcd[15:4]};

//������ʾʹ�ܣ���λ����
assign dat_en[7] = |T_data[15:12]; //�Ի�
assign dat_en[6] = (b>=32'd4685)?(|T_data[15:8]):(|T_data[11:8]);
assign dat_en[5:4] = 2'b11;

//С������ʾʹ��
assign dot_en[7:4] = 4'b0010;

/////////////////////////////////////ʪ������/////////////////////////////////////////

// ʪ�� TH = -6 + 125 * H_code / 2^16 = (-60 + 1250 * H_code / 2^16) / 10
wire [31:0] d = H_code * 16'd1250;
wire [31:0] e = d >> 16; //����2^16ȡ��
wire [31:0] f = e - 32'd60;
wire [15:0] H_data_bin = f[15:0];

//����BCDת�봦��
//С������BCD�����������1λ����ɳ���10�Ĳ���
//H_data_bcd[19:16]ǧλ,[15:12]��λ,[11:8]ʮλ,[7:4]��λ,[3:0]С��λ
wire [19:0] H_data_bcd;
bin_to_bcd u2
(
.rst_n				(rst_n		),	//ϵͳ��λ������Ч
.bin_code			(H_data_bin	),	//��Ҫ����BCDת��Ķ���������
.bcd_code			(H_data_bcd	)	//ת����BCD�����������
);

//Ҫ��ʾ������,����1λС��
assign H_data = H_data_bcd[15:0];

//������ʾʹ��
assign dat_en[3] = |H_data[15:12]; //�Ի�
assign dat_en[2] = |H_data[15:8];
assign dat_en[1:0] = 2'b11;

//С������ʾʹ��
assign dot_en[3:0] = 4'b0010;

endmodule
