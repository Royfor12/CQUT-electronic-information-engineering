// ********************************************************************
// >>>>>>>>>>>>>>>>>>>>>>>>> COPYRIGHT NOTICE <<<<<<<<<<<<<<<<<<<<<<<<<
// ********************************************************************
// File name    : decode38.v
// Module name  : decode38
// Author       : STEP
// Description  : 3-8decode control LED
// Web          : www.stepfpga.com
// 
// --------------------------------------------------------------------
// Code Revision History : 
// --------------------------------------------------------------------
// Version: |Mod. Date:   |Changes Made:
// V1.0     |2017/03/02   |Initial ver
// --------------------------------------------------------------------
// Module Function:����3·���ص�״̬��Ϊ�����ͨ��3-8����ʵ�ֿ���LED�Ƶ���ʾ��
 
module decode38 (sw,led);
 
	input [2:0] sw;		//���������źţ�����������3��������Ϊ3-8������������
	output [7:0] led;	//����źſ����ض�LED
 
        reg [7:0] led;  //����ledΪreg�ͱ�������always���̿���ֻ�ܶ�reg�ͱ�����ֵ
 
    //always���̿飬������swΪ���б�������sw�仯һ��ִ��һ��always��������䣬���򱣳ֲ���
	always @ (sw)
	begin
		case(sw)                       //case��䣬һ��Ҫ��default���
			3'b000:	led=8'b0111_1111;  //������ת�����С�_���»���ֻ��Ϊ���Ķ����㣬��ʵ������  
			3'b001:	led=8'b1011_1111;  //λ��'����+��ֵ��Verilog�ﳣ���ı�﷽�������ƿ�����b��o��d��h�������ˡ�ʮ��ʮ�����ƣ�
			3'b010:	led=8'b1101_1111;
			3'b011:	led=8'b1110_1111;
			3'b100:	led=8'b1111_0111;
			3'b101:	led=8'b1111_1011;
			3'b110: led=8'b1111_1101;
			3'b111:	led=8'b1111_1110;
			default: ;
		endcase
	end
 
endmodule